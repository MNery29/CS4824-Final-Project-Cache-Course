// Test Module for rob unit


`include "verilog/sys_defs.svh"