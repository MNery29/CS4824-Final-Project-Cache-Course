// tests to do:
