// dummy for testing