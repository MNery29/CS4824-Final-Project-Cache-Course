/*
dcache specifications:
    256-bytes, 32 lines
    non-blocking
    write-back
    set-associative
    z-cache design -- https://people.csail.mit.edu/sanchez/papers/2010.zcache.micro.pdf

*/