// Test Module for rob unit


`include "verilog/sys_defs.svh"

// Tests to include: 

// Test for full capacity of the ROB
